`define OP_LOAD 4'd0
`define OP_SHIFT_R 4'd1
`define OP_SHIFT_L 4'd2
`define OP_SHIFT_U 4'd3
`define OP_SHIFT_D 4'd4
`define OP_REDUCE 4'd5
`define OP_INCREASE 4'd6
`define OP_DISPLAY 4'd7
`define OP_CONV 4'd8
`define OP_MEDIAN 4'd9
`define OP_SGNMS 4'd10
`define ORIGIN_COL origin[2:0]
`define ORIGIN_ROW origin[5:3] 
`define PE_CONV1_4 4'd0
`define PE_CONV1_8 4'd1
`define PE_CONV1_16 4'd2
`define PE_NMS2 4'd3
`define PE_NMS1 4'd4
`define PE_NMS0 4'd5
`define PE_NMS_1 4'd6
`define PE_NMS_2 4'd7
`define PE_MED 4'd8
`define ANGLE0 2'd0
`define ANGLE45 2'd1
`define ANGLE90 2'd2
`define ANGLE135 2'd3